 -- constant here : audio_incnv_t := 2+3;  -- use in clear statements
 -- constant there : audio_incnv_t := 2+5;  
  constant oops : audio_incnv_t := "01111011";  