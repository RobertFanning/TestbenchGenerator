package ${NAME}_type_pkg;
Fetch_Interface:
IncludePackages:
//DEFINE UNPACKED TYPES AS SYSTEMVERILOG FORMAT
Type_Package_Unpacked:

//DEFINE VIRTUAL INTERFACE TYPES HERE
Fetch_Interface:
type_pkg_virtual_interface:


endpackage;
