constant C_SCALING_VEC_LEN : positive := 3;
subtype scaling_t is unsigned(C_SCALING_VEC_LEN-1 downto 0)