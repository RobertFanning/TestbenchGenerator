constant C_X_DECODED_ZERO : x_decoded_t := 1+2*3;
